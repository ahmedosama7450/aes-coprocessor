module tb_aes;
    tb_wrapper #(.WITH_AES(1'b1)) tb ();
endmodule
