module tb;
    tb_wrapper #(.WITH_AES(1'b0)) tb ();
endmodule
